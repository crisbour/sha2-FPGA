`define CODEC_POS            32     // Tuser position: 32nd bit in tuser in begining of user_slot_0 taken by codec

// Used define codecs
`define CODEC_SHA2_224        16'h09
`define CODEC_SHA2_384        16'h10

// Hash codecs
`define CODEC_SHA1            16'h11
`define CODEC_SHA2_256        16'h12
`define CODEC_SHA2_512        16'h13
`define CODEC_SHA3_512        16'h14
`define CODEC_SHA3_384        16'h15
`define CODEC_SHA3_256        16'h16
`define CODEC_SHA3_224        16'h17
`define CODEC_SHAKE_128       16'h18
`define CODEC_SHAKE_256       16'h19
`define CODEC_KECCAK_224      16'h1A
`define CODEC_KECCAK_256      16'h1B
`define CODEC_KECCAK_384      16'h1C
`define CODEC_KECCAK_512      16'h1D
`define CODEC_BLAKE3          16'h1E
`define CODEC_DCCP            16'h21
`define CODEC_MURMUR3_128     16'h22
`define CODEC_DBL_SHA2_256    16'h56
`define CODEC_MD4             16'hD4
`define CODEC_MD5             16'hD5
`define CODEC_BMT             16'hD6
`define CODEC_SHA2_256_TRUNC254_PADDED      16'h1012
`define CODEC_RIPEMD_128      16'h1052
`define CODEC_RIPEMD_160      16'h1053
`define CODEC_RIPEMD_256      16'h1054
`define CODEC_RIPEMD_320      16'h1055
`define CODEC_X11             16'h1100
`define CODEC_KANGAROOTWELVE  16'h1D01
`define CODEC_SM3_256         16'h534D
`define CODEC_BLAKE2B_8       16'hB201
`define CODEC_BLAKE2B_16      16'hB202
`define CODEC_BLAKE2B_24      16'hB203
`define CODEC_BLAKE2B_32      16'hB204
`define CODEC_BLAKE2B_40      16'hB205
`define CODEC_BLAKE2B_48      16'hB206
`define CODEC_BLAKE2B_56      16'hB207
`define CODEC_BLAKE2B_64      16'hB208
`define CODEC_BLAKE2B_72      16'hB209
`define CODEC_BLAKE2B_80      16'hB20A
`define CODEC_BLAKE2B_88      16'hB20B
`define CODEC_BLAKE2B_96      16'hB20C
`define CODEC_BLAKE2B_104      16'hB20D
`define CODEC_BLAKE2B_112      16'hB20E
`define CODEC_BLAKE2B_120      16'hB20F
`define CODEC_BLAKE2B_128      16'hB210
`define CODEC_BLAKE2B_136      16'hB211
`define CODEC_BLAKE2B_144      16'hB212
`define CODEC_BLAKE2B_152      16'hB213
`define CODEC_BLAKE2B_160      16'hB214
`define CODEC_BLAKE2B_168      16'hB215
`define CODEC_BLAKE2B_176      16'hB216
`define CODEC_BLAKE2B_184      16'hB217
`define CODEC_BLAKE2B_192      16'hB218
`define CODEC_BLAKE2B_200      16'hB219
`define CODEC_BLAKE2B_208      16'hB21A
`define CODEC_BLAKE2B_216      16'hB21B
`define CODEC_BLAKE2B_224      16'hB21C
`define CODEC_BLAKE2B_232      16'hB21D
`define CODEC_BLAKE2B_240      16'hB21E
`define CODEC_BLAKE2B_248      16'hB21F
`define CODEC_BLAKE2B_256      16'hB220
`define CODEC_BLAKE2B_264      16'hB221
`define CODEC_BLAKE2B_272      16'hB222
`define CODEC_BLAKE2B_280      16'hB223
`define CODEC_BLAKE2B_288      16'hB224
`define CODEC_BLAKE2B_296      16'hB225
`define CODEC_BLAKE2B_304      16'hB226
`define CODEC_BLAKE2B_312      16'hB227
`define CODEC_BLAKE2B_320      16'hB228
`define CODEC_BLAKE2B_328      16'hB229
`define CODEC_BLAKE2B_336      16'hB22A
`define CODEC_BLAKE2B_344      16'hB22B
`define CODEC_BLAKE2B_352      16'hB22C
`define CODEC_BLAKE2B_360      16'hB22D
`define CODEC_BLAKE2B_368      16'hB22E
`define CODEC_BLAKE2B_376      16'hB22F
`define CODEC_BLAKE2B_384      16'hB230
`define CODEC_BLAKE2B_392      16'hB231
`define CODEC_BLAKE2B_400      16'hB232
`define CODEC_BLAKE2B_408      16'hB233
`define CODEC_BLAKE2B_416      16'hB234
`define CODEC_BLAKE2B_424      16'hB235
`define CODEC_BLAKE2B_432      16'hB236
`define CODEC_BLAKE2B_440      16'hB237
`define CODEC_BLAKE2B_448      16'hB238
`define CODEC_BLAKE2B_456      16'hB239
`define CODEC_BLAKE2B_464      16'hB23A
`define CODEC_BLAKE2B_472      16'hB23B
`define CODEC_BLAKE2B_480      16'hB23C
`define CODEC_BLAKE2B_488      16'hB23D
`define CODEC_BLAKE2B_496      16'hB23E
`define CODEC_BLAKE2B_504      16'hB23F
`define CODEC_BLAKE2B_512      16'hB240
`define CODEC_BLAKE2S_8       16'hB241
`define CODEC_BLAKE2S_16      16'hB242
`define CODEC_BLAKE2S_24      16'hB243
`define CODEC_BLAKE2S_32      16'hB244
`define CODEC_BLAKE2S_40      16'hB245
`define CODEC_BLAKE2S_48      16'hB246
`define CODEC_BLAKE2S_56      16'hB247
`define CODEC_BLAKE2S_64      16'hB248
`define CODEC_BLAKE2S_72      16'hB249
`define CODEC_BLAKE2S_80      16'hB24A
`define CODEC_BLAKE2S_88      16'hB24B
`define CODEC_BLAKE2S_96      16'hB24C
`define CODEC_BLAKE2S_104      16'hB24D
`define CODEC_BLAKE2S_112      16'hB24E
`define CODEC_BLAKE2S_120      16'hB24F
`define CODEC_BLAKE2S_128      16'hB250
`define CODEC_BLAKE2S_136      16'hB251
`define CODEC_BLAKE2S_144      16'hB252
`define CODEC_BLAKE2S_152      16'hB253
`define CODEC_BLAKE2S_160      16'hB254
`define CODEC_BLAKE2S_168      16'hB255
`define CODEC_BLAKE2S_176      16'hB256
`define CODEC_BLAKE2S_184      16'hB257
`define CODEC_BLAKE2S_192      16'hB258
`define CODEC_BLAKE2S_200      16'hB259
`define CODEC_BLAKE2S_208      16'hB25A
`define CODEC_BLAKE2S_216      16'hB25B
`define CODEC_BLAKE2S_224      16'hB25C
`define CODEC_BLAKE2S_232      16'hB25D
`define CODEC_BLAKE2S_240      16'hB25E
`define CODEC_BLAKE2S_248      16'hB25F
`define CODEC_BLAKE2S_256      16'hB260
`define CODEC_SKEIN256_8       16'hB301
`define CODEC_SKEIN256_16      16'hB302
`define CODEC_SKEIN256_24      16'hB303
`define CODEC_SKEIN256_32      16'hB304
`define CODEC_SKEIN256_40      16'hB305
`define CODEC_SKEIN256_48      16'hB306
`define CODEC_SKEIN256_56      16'hB307
`define CODEC_SKEIN256_64      16'hB308
`define CODEC_SKEIN256_72      16'hB309
`define CODEC_SKEIN256_80      16'hB30A
`define CODEC_SKEIN256_88      16'hB30B
`define CODEC_SKEIN256_96      16'hB30C
`define CODEC_SKEIN256_104      16'hB30D
`define CODEC_SKEIN256_112      16'hB30E
`define CODEC_SKEIN256_120      16'hB30F
`define CODEC_SKEIN256_128      16'hB310
`define CODEC_SKEIN256_136      16'hB311
`define CODEC_SKEIN256_144      16'hB312
`define CODEC_SKEIN256_152      16'hB313
`define CODEC_SKEIN256_160      16'hB314
`define CODEC_SKEIN256_168      16'hB315
`define CODEC_SKEIN256_176      16'hB316
`define CODEC_SKEIN256_184      16'hB317
`define CODEC_SKEIN256_192      16'hB318
`define CODEC_SKEIN256_200      16'hB319
`define CODEC_SKEIN256_208      16'hB31A
`define CODEC_SKEIN256_216      16'hB31B
`define CODEC_SKEIN256_224      16'hB31C
`define CODEC_SKEIN256_232      16'hB31D
`define CODEC_SKEIN256_240      16'hB31E
`define CODEC_SKEIN256_248      16'hB31F
`define CODEC_SKEIN256_256      16'hB320
`define CODEC_SKEIN512_8       16'hB321
`define CODEC_SKEIN512_16      16'hB322
`define CODEC_SKEIN512_24      16'hB323
`define CODEC_SKEIN512_32      16'hB324
`define CODEC_SKEIN512_40      16'hB325
`define CODEC_SKEIN512_48      16'hB326
`define CODEC_SKEIN512_56      16'hB327
`define CODEC_SKEIN512_64      16'hB328
`define CODEC_SKEIN512_72      16'hB329
`define CODEC_SKEIN512_80      16'hB32A
`define CODEC_SKEIN512_88      16'hB32B
`define CODEC_SKEIN512_96      16'hB32C
`define CODEC_SKEIN512_104      16'hB32D
`define CODEC_SKEIN512_112      16'hB32E
`define CODEC_SKEIN512_120      16'hB32F
`define CODEC_SKEIN512_128      16'hB330
`define CODEC_SKEIN512_136      16'hB331
`define CODEC_SKEIN512_144      16'hB332
`define CODEC_SKEIN512_152      16'hB333
`define CODEC_SKEIN512_160      16'hB334
`define CODEC_SKEIN512_168      16'hB335
`define CODEC_SKEIN512_176      16'hB336
`define CODEC_SKEIN512_184      16'hB337
`define CODEC_SKEIN512_192      16'hB338
`define CODEC_SKEIN512_200      16'hB339
`define CODEC_SKEIN512_208      16'hB33A
`define CODEC_SKEIN512_216      16'hB33B
`define CODEC_SKEIN512_224      16'hB33C
`define CODEC_SKEIN512_232      16'hB33D
`define CODEC_SKEIN512_240      16'hB33E
`define CODEC_SKEIN512_248      16'hB33F
`define CODEC_SKEIN512_256      16'hB340
`define CODEC_SKEIN512_264      16'hB341
`define CODEC_SKEIN512_272      16'hB342
`define CODEC_SKEIN512_280      16'hB343
`define CODEC_SKEIN512_288      16'hB344
`define CODEC_SKEIN512_296      16'hB345
`define CODEC_SKEIN512_304      16'hB346
`define CODEC_SKEIN512_312      16'hB347
`define CODEC_SKEIN512_320      16'hB348
`define CODEC_SKEIN512_328      16'hB349
`define CODEC_SKEIN512_336      16'hB34A
`define CODEC_SKEIN512_344      16'hB34B
`define CODEC_SKEIN512_352      16'hB34C
`define CODEC_SKEIN512_360      16'hB34D
`define CODEC_SKEIN512_368      16'hB34E
`define CODEC_SKEIN512_376      16'hB34F
`define CODEC_SKEIN512_384      16'hB350
`define CODEC_SKEIN512_392      16'hB351
`define CODEC_SKEIN512_400      16'hB352
`define CODEC_SKEIN512_408      16'hB353
`define CODEC_SKEIN512_416      16'hB354
`define CODEC_SKEIN512_424      16'hB355
`define CODEC_SKEIN512_432      16'hB356
`define CODEC_SKEIN512_440      16'hB357
`define CODEC_SKEIN512_448      16'hB358
`define CODEC_SKEIN512_456      16'hB359
`define CODEC_SKEIN512_464      16'hB35A
`define CODEC_SKEIN512_472      16'hB35B
`define CODEC_SKEIN512_480      16'hB35C
`define CODEC_SKEIN512_488      16'hB35D
`define CODEC_SKEIN512_496      16'hB35E
`define CODEC_SKEIN512_504      16'hB35F
`define CODEC_SKEIN512_512      16'hB360
`define CODEC_SKEIN1024_8       16'hB361
`define CODEC_SKEIN1024_16      16'hB362
`define CODEC_SKEIN1024_24      16'hB363
`define CODEC_SKEIN1024_32      16'hB364
`define CODEC_SKEIN1024_40      16'hB365
`define CODEC_SKEIN1024_48      16'hB366
`define CODEC_SKEIN1024_56      16'hB367
`define CODEC_SKEIN1024_64      16'hB368
`define CODEC_SKEIN1024_72      16'hB369
`define CODEC_SKEIN1024_80      16'hB36A
`define CODEC_SKEIN1024_88      16'hB36B
`define CODEC_SKEIN1024_96      16'hB36C
`define CODEC_SKEIN1024_104      16'hB36D
`define CODEC_SKEIN1024_112      16'hB36E
`define CODEC_SKEIN1024_120      16'hB36F
`define CODEC_SKEIN1024_128      16'hB370
`define CODEC_SKEIN1024_136      16'hB371
`define CODEC_SKEIN1024_144      16'hB372
`define CODEC_SKEIN1024_152      16'hB373
`define CODEC_SKEIN1024_160      16'hB374
`define CODEC_SKEIN1024_168      16'hB375
`define CODEC_SKEIN1024_176      16'hB376
`define CODEC_SKEIN1024_184      16'hB377
`define CODEC_SKEIN1024_192      16'hB378
`define CODEC_SKEIN1024_200      16'hB379
`define CODEC_SKEIN1024_208      16'hB37A
`define CODEC_SKEIN1024_216      16'hB37B
`define CODEC_SKEIN1024_224      16'hB37C
`define CODEC_SKEIN1024_232      16'hB37D
`define CODEC_SKEIN1024_240      16'hB37E
`define CODEC_SKEIN1024_248      16'hB37F
`define CODEC_SKEIN1024_256      16'hB380
`define CODEC_SKEIN1024_264      16'hB381
`define CODEC_SKEIN1024_272      16'hB382
`define CODEC_SKEIN1024_280      16'hB383
`define CODEC_SKEIN1024_288      16'hB384
`define CODEC_SKEIN1024_296      16'hB385
`define CODEC_SKEIN1024_304      16'hB386
`define CODEC_SKEIN1024_312      16'hB387
`define CODEC_SKEIN1024_320      16'hB388
`define CODEC_SKEIN1024_328      16'hB389
`define CODEC_SKEIN1024_336      16'hB38A
`define CODEC_SKEIN1024_344      16'hB38B
`define CODEC_SKEIN1024_352      16'hB38C
`define CODEC_SKEIN1024_360      16'hB38D
`define CODEC_SKEIN1024_368      16'hB38E
`define CODEC_SKEIN1024_376      16'hB38F
`define CODEC_SKEIN1024_384      16'hB390
`define CODEC_SKEIN1024_392      16'hB391
`define CODEC_SKEIN1024_400      16'hB392
`define CODEC_SKEIN1024_408      16'hB393
`define CODEC_SKEIN1024_416      16'hB394
`define CODEC_SKEIN1024_424      16'hB395
`define CODEC_SKEIN1024_432      16'hB396
`define CODEC_SKEIN1024_440      16'hB397
`define CODEC_SKEIN1024_448      16'hB398
`define CODEC_SKEIN1024_456      16'hB399
`define CODEC_SKEIN1024_464      16'hB39A
`define CODEC_SKEIN1024_472      16'hB39B
`define CODEC_SKEIN1024_480      16'hB39C
`define CODEC_SKEIN1024_488      16'hB39D
`define CODEC_SKEIN1024_496      16'hB39E
`define CODEC_SKEIN1024_504      16'hB39F
`define CODEC_SKEIN1024_512      16'hB3A0
`define CODEC_SKEIN1024_520      16'hB3A1
`define CODEC_SKEIN1024_528      16'hB3A2
`define CODEC_SKEIN1024_536      16'hB3A3
`define CODEC_SKEIN1024_544      16'hB3A4
`define CODEC_SKEIN1024_552      16'hB3A5
`define CODEC_SKEIN1024_560      16'hB3A6
`define CODEC_SKEIN1024_568      16'hB3A7
`define CODEC_SKEIN1024_576      16'hB3A8
`define CODEC_SKEIN1024_584      16'hB3A9
`define CODEC_SKEIN1024_592      16'hB3AA
`define CODEC_SKEIN1024_600      16'hB3AB
`define CODEC_SKEIN1024_608      16'hB3AC
`define CODEC_SKEIN1024_616      16'hB3AD
`define CODEC_SKEIN1024_624      16'hB3AE
`define CODEC_SKEIN1024_632      16'hB3AF
`define CODEC_SKEIN1024_640      16'hB3B0
`define CODEC_SKEIN1024_648      16'hB3B1
`define CODEC_SKEIN1024_656      16'hB3B2
`define CODEC_SKEIN1024_664      16'hB3B3
`define CODEC_SKEIN1024_672      16'hB3B4
`define CODEC_SKEIN1024_680      16'hB3B5
`define CODEC_SKEIN1024_688      16'hB3B6
`define CODEC_SKEIN1024_696      16'hB3B7
`define CODEC_SKEIN1024_704      16'hB3B8
`define CODEC_SKEIN1024_712      16'hB3B9
`define CODEC_SKEIN1024_720      16'hB3BA
`define CODEC_SKEIN1024_728      16'hB3BB
`define CODEC_SKEIN1024_736      16'hB3BC
`define CODEC_SKEIN1024_744      16'hB3BD
`define CODEC_SKEIN1024_752      16'hB3BE
`define CODEC_SKEIN1024_760      16'hB3BF
`define CODEC_SKEIN1024_768      16'hB3C0
`define CODEC_SKEIN1024_776      16'hB3C1
`define CODEC_SKEIN1024_784      16'hB3C2
`define CODEC_SKEIN1024_792      16'hB3C3
`define CODEC_SKEIN1024_800      16'hB3C4
`define CODEC_SKEIN1024_808      16'hB3C5
`define CODEC_SKEIN1024_816      16'hB3C6
`define CODEC_SKEIN1024_824      16'hB3C7
`define CODEC_SKEIN1024_832      16'hB3C8
`define CODEC_SKEIN1024_840      16'hB3C9
`define CODEC_SKEIN1024_848      16'hB3CA
`define CODEC_SKEIN1024_856      16'hB3CB
`define CODEC_SKEIN1024_864      16'hB3CC
`define CODEC_SKEIN1024_872      16'hB3CD
`define CODEC_SKEIN1024_880      16'hB3CE
`define CODEC_SKEIN1024_888      16'hB3CF
`define CODEC_SKEIN1024_896      16'hB3D0
`define CODEC_SKEIN1024_904      16'hB3D1
`define CODEC_SKEIN1024_912      16'hB3D2
`define CODEC_SKEIN1024_920      16'hB3D3
`define CODEC_SKEIN1024_928      16'hB3D4
`define CODEC_SKEIN1024_936      16'hB3D5
`define CODEC_SKEIN1024_944      16'hB3D6
`define CODEC_SKEIN1024_952      16'hB3D7
`define CODEC_SKEIN1024_960      16'hB3D8
`define CODEC_SKEIN1024_968      16'hB3D9
`define CODEC_SKEIN1024_976      16'hB3DA
`define CODEC_SKEIN1024_984      16'hB3DB
`define CODEC_SKEIN1024_992      16'hB3DC
`define CODEC_SKEIN1024_1000      16'hB3DD
`define CODEC_SKEIN1024_1008      16'hB3DE
`define CODEC_SKEIN1024_1016      16'hB3DF
`define CODEC_SKEIN1024_1024      16'hB3E0
`define CODEC_POSEIDON_BLS12_381_A2_FC1         16'hB401
`define CODEC_POSEIDON_BLS12_381_A2_FC1_SC      16'hB402

// Multihash codec
`define CODEC_MULTIHASH       16'h31
